module adder_pc(input[31:0] operando_1, input[31:0] operando_2, output [31:0] resultado);

assing y = operando_1 + operando_2;

endmodule
	