library verilog;
use verilog.vl_types.all;
entity tb_extensor is
end tb_extensor;
