library verilog;
use verilog.vl_types.all;
entity tb_cont_prog is
end tb_cont_prog;
