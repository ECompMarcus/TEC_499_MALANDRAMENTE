library verilog;
use verilog.vl_types.all;
entity tb_memoria is
end tb_memoria;
