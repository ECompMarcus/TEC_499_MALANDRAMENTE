`ifndef ALUOP
`define ALUOP

`define ALU_ADDU 5'd0
`define ALU_SUBU 5'd1
`define ALU_SLT  5'd2
`define ALU_SLTU 5'd3
`define ALU_AND  5'd4
`define ALU_OR   5'd5
`define ALU_XOR  5'd6
`define ALU_LUI  5'd7
`define ALU_SLL  5'd8
`define ALU_SRL  5'd9
`define ALU_SRA  5'd10
`define ALU_NOR  5'd11
//ADCIONADAS
`define ALU_SUB	5'd12
`define ALU_ADD	5'd13
//`define ALU_SLA 	5'd14
`define ALU_BEQ  	5'd15
`define ALU_BNE  	5'd16
`define ALU_BLEZ  5'd17
`define ALU_BGTZ  5'd18
`define ALU_BLTZ  5'd19
`define ALU_BGEZ  5'd20
`define ALU_CLZ  	5'd21
`define ALU_CLO  	5'd22

`define ALU_XXX  5'd26

`endif //ALUOP
