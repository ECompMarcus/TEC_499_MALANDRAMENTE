library verilog;
use verilog.vl_types.all;
entity tb_banco is
end tb_banco;
